/*#############################################################################\
##                                                                            ##
##       Applied Electronics - Physics Department - University of Padova      ##
##                                                                            ##
\#############################################################################*/

// Set timescale (default time unit if not otherwise specified).
`timescale 1ns / 1ps

// Emulate a DS ADC
module adc_emulator (
    input CLK,
    input RST_B,
    output DRIVE
    );
endmodule
